ARCHITECTURE masterVersion OF offsetAdd IS
BEGIN
  phaseOut <= offset + phaseIn;
END ARCHITECTURE masterVersion;
